* Лабораторная работа №2
* ----------------------
* Симметричный мультивибратор с нагрузкой на светодиоды

* источник питания +4.5В
VCC VCC 0 DC 4.5V

* конденсаторы
C1 vc1 vb2 22uF  
C2 vc2 vb1 22uF  

* резисторы
R1 vc1 VCC 1k  
R2 vb2 VCC 33k  
R3 vb1 VCC 33k  
R4 vc2 VCC 1k  
R5 vc3 vled1 57  
R6 vc4 vled2 57  

* транзисторы
QVT1 vc1 vb1 ve1 2N2222 
QVT2 vc2 vb2 ve2 2N2222 
QVT3 vc3 ve1 0 2N2222 
QVT4 vc4 ve2 0 2N2222 

* светодиоды
DLED1 VCC vled1 NSPW500BS 
DLED2 VCC vled2 NSPW500BS 

* SPICE модель классического импортного транзистора 2N2222
.model 2N2222 NPN (IS=19.34n EG=1.11 VAF=250.3 BF=163.8 ISE =174.3f
+  NE=1.647 IKF=3.0 XTB=1.5 BR=11.49 ISC=19.9f NC=1.88 IKR=10.75
+  RC=0.3567 CJC=11.02p VJC=0.3869 MJC=0.3292 FC=0.5 CJE=29.31p VJE=0.9036
+  MJE=0.4101 TR=38.32n TF=361.8p ITF=5.282 XTF=249.9 VTF=10)

* SPICE модель "стандартного" светодиода NSPW500BS
.model NSPW500BS D(Is=.27n Rs=5.65 N=6.79 Cjo=42p Xti=200)

* температурный режим
.options TEMP=25

* моделирование переходного процесса
* шаг моделирования - 1 мс
* время моделирования - 10 с
.tran 1m 10

.end

