* File: "lab-4.cir"
* Работа биполярного транзистора в нелинейном (импульсном) режиме.

* источник питания +5В
VCC vcc 0 DC 5V

* источник сигнала
VSIN vpulse 0 dc 0V ac 1mV pulse(0V 2V 0.4ms 0.1ms 0.1ms 0.33ms 1ms)

* внутреннее сопротивление источника сигнала
RIN vpulse vin 75

* входной конденсатор
CIN vin vcin 10uF

* импульсный диод для восстановления постоянной составляющей
D1 0 vcin 1N914
*R2 0 vcin 1k

* резистор - ограничитель тока базы
RB vcin vbb 220

* фиктивный источик напряжения 0В для контроля базового тока
VB vbb vb 0V

* n-p-n транзистор
QT1 vc vb 0 2T325V

* фиктивный источик напряжения 0В для контроля базового тока
VC vc vvc 0V

* резистор-нагрузка к коллекторной цепи транзистора
RL vcc vvc 1k

* SPICE модель советского "военного" транзистора 2T325В (h21э=321.5) 
.model 2T325V NPN(Is=9.164f Xti=3 Eg=1.11 Vaf=87 Bf=321.5 Ise=87.74f 
+  Ne=1.473 Ikf=87.77m Xtb=1.5 Br=1.78 Isc=.1p Nc=1.744 Ikr=.6068
+  Rb=31 Rc=.2997 Cjc=2.958p Mjc=.333 Vjc=.75 Fc=.5 Cje=3.42p Mje=.333
+  Vje=.75 Tr=8.891n Tf=112.2p Itf=.3 Xtf=2 Vtf=25)

* SPICE модель кремневого диода 1N914/1N4148 - аналог КД521А
.model 1N914 D(Is=2.52n Rs=.568 N=1.752 Cjo=4p M=.4 tt=20n)

* температурный режим
.options TEMP=27

* моделирование переходного процесса
* шаг моделирования - 1 мкс
* время моделирования - 30 мс
.tran 1u 30m

.end

