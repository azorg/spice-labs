* Лабораторная работа №3
* ----------------------
* Измерение входных и выходных вольт-амперных характеристик (ВАХ)
* SPICE модели биполярного транзистора

* напряжение на коллекторе (0..15В)
VC vc 0 DC 5V

* напряжение на базе (при снятии входной ВАХ)
VB vb 0 DC 0.5V

* ИЛИ

* ток базы (при снятии выходной ВАХ и при снятии зависимости Ic(Ib))
*IB 0 vb DC 1uA

* NPN транзистор
QVT vc vb 0 KT315B

* SPICE модель классического советского транзистора КТ315Б (h21э~100)
.model KT315B NPN(Is=14.34f Xti=3 Eg=1.11 Vaf=125 Bf=124 Ise=157.3f
+  Ne=1.558 Ikf=.2999 Xtb=1.5 Br=1 Isc=15.86f Nc=1.022
+  Ikr=3.163 Rb=15 Rc=3.748 Cjc=8.988p Mjc=.33 Vjc=.75 Fc=.5 Cje=18.5p
+  Mje=.33 Vje=.75 Tr=301.4n Tf=321.4p Itf=1 Xtf=2 Vtf=60)

* температурный режим
.options TEMP=25

.end

