* File: "lab-11.cir"
* Несимметричный мультивибратор - генератор коротких импульсов

* источник питания +4.5В
VCC VCC 0 DC 4.5V

* конденсатор
C1 v1 vc2 22uF

* резисторы
R1 VCC  v1   68k
R2 vb1  v1   1k
R3 vb1  0    10k
R4 vc1  vb2  10k  
R5 vc2  0    2.2k
R6 vc2  vled 150

* транзисторы
QVT1 vc1 vb1 0   2N3904
QVT2 vc2 vb2 VCC 2N3906

* светодиод
DLED1 vled 0 NSPW500BS 

* SPICE модель транзистора 2N3904 (из просторов Интернет):
.MODEL 2N3904 npn
+IS=6.9716e-14 BF=545.416 NF=1.09328 VAF=10
+IKF=0.0228393 ISE=5.71808e-12 NE=1.88204 BR=4.70256
+NR=1.3912 VAR=2.31769 IKR=0.074093 ISC=5.71808e-12
+NC=1.36259 RB=1.733 IRB=1.12054 RBM=0.876202
+RE=0.356192 RC=1.78096 XTB=0.1 XTI=1
+EG=1.05 CJE=4.47982e-12 VJE=0.4 MJE=0.240345
+TF=4e-10 XTF=1.5 VTF=1 ITF=1
+CJC=3.76637e-12 VJC=0.4 MJC=0.241382 XCJC=0.8
+FC=0.533333 CJS=0 VJS=0.75 MJS=0.5
+TR=3.77901e-05 PTF=0 KF=0 AF=1

* SPICE модель транзистора 2N3906 (из просторов Интернет):
.MODEL 2N3906 PNP
+IS=1.14615e-14 BF=535.453 NF=1.06473 VAF=10
+IKF=0.0234918 ISE=1.33613e-13 NE=1.62939 BR=4.66099
+NR=1.19618 VAR=2.77165 IKR=0.0740931 ISC=1.33613e-13
+NC=1.22182 RB=0.1 IRB=1.05964 RBM=0.1
+RE=0.0001 RC=1.39183 XTB=0.1 XTI=1
+EG=1.05 CJE=6.03788e-12 VJE=0.4 MJE=0.272764
+TF=4.8381e-10 XTF=1.5 VTF=1 ITF=1
+CJC=6.18444e-12 VJC=0.4 MJC=0.234098 XCJC=0.8
+FC=0.5415 CJS=0 VJS=0.75 MJS=0.5
+TR=2.42096e-06 PTF=0 KF=0 AF=1

* SPICE модель "стандартного" светодиода NSPW500BS
.model NSPW500BS D(Is=.27n Rs=5.65 N=6.79 Cjo=42p Xti=200)

* температурный режим
.options TEMP=25

* моделирование переходного процесса
* шаг моделирования - 50 мкс
* время моделирования - 5 с
.tran 50u 5

.end

