* File: "lab-1.cir"
* Усилитель переменного тока на 2-х биполярных транзисторах с непосредственными
* связями по схеме ОЭ и ОК с обратной отрицательной связью по постоянному
* и переменному току.

* конденсаторы
CIN vin vb 10uF  
COUT ve2 vout 100uF
CE 0 vce 33uF  
CCOR ve vce 10pF
CVCC VCC 0 1000uF  

* дроссель частотной коррекции в коллекторной цепи VT1
LCOR vl vc 33uH

* резисторы
R1 vb VCC 30k
R2 0 vb 10k
R3 vl VCC 3.3k
R4 ve vce 200
R5 0 vce 1k
R6 0 ve2 470

* внутреннее сопротивление источника
RIN vsin vin 1k

* сопротивление нагрузки
RL 0 vout 1000

* источник питания +9В
VCC vcc 0 DC 9V

* источник сигнала
VSIN vsin 0 dc 0 ac 1mV sin(0 1mV 1kHz)

* n-p-n транзисторы
QVT1 vc  vb ve  KT368B
QVT2 VCC vc ve2 KT368B

* SPICE модель советского ВЧ транзистора КТ368Б (h21э=110)
.model KT368B NPN(Is=8.675f Xti=3 Eg=1.11 Vaf=108 Bf=110 Ne=1.377
+  Ise=9.128f Ikf=.3608 Xtb=1.5 Var=56 Br=1.45 Nc=2 Isc=16.3f Ikr=.125
+  Rb=31.5 Rc=2.445 Cjc=2.35p Vjc=.75 Mjc=.33 Fc=.5 Cje=2.786p Vje=.69
+  Mje=.37 Tr=2.147n Tf=84.62p Itf=.15 Vtf=25 Xtf=2)

* температурный режим
.options TEMP=25

* моделирование переходного процесса
* шаг моделирования - 1 мкс
* время моделирования - 10 мс
.tran 1u 10m

.end

