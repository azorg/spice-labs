* File: "lab-3_2.cir"
* Измерение выходных вольт-амперных характеристик (ВАХ) 
* SPICE модели биполярного транзистора

* токи баз транзисторов
IB1 0 vb1 DC 10uA
IB2 0 vb2 DC 50uA
IB3 0 vb3 DC 100uA

* напряжение на коллекторах транзисторов
VC vc 0 DC 5V

* фиктивные источники нулевого напряжения для измерения токов коллекторов
VC1 vc vc1 DC 0V
VC2 vc vc2 DC 0V
VC3 vc vc3 DC 0V

* идентичные n-p-n транзисторы с разными токами базы
QVT1 vc1 vb1 0 KT315B
QVT2 vc2 vb2 0 KT315B
QVT3 vc3 vb3 0 KT315B

* SPICE модель классического советского транзистора КТ315Б (h21э=100)
.model KT315B NPN(Is=14.34f Xti=3 Eg=1.11 Vaf=125 Bf=124 Ise=157.3f
+  Ne=1.558 Ikf=.2999 Xtb=1.5 Br=1 Isc=15.86f Nc=1.022
+  Ikr=3.163 Rb=15 Rc=3.748 Cjc=8.988p Mjc=.33 Vjc=.75 Fc=.5 Cje=18.5p
+  Mje=.33 Vje=.75 Tr=301.4n Tf=321.4p Itf=1 Xtf=2 Vtf=60)

* температурный режим
.options TEMP=27

* DC анализ при различном напряжении на коллекторах (0...15В)
.dc vc 0V 15V 1mV

* Графики зависимости тока коллектора от напряжения на коллекторе
* -> run
* -> plot i(vc1) i(vc2) i(vc3)

.end

