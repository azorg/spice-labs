* File: "sandbox.cir"
* Простые схемы для проверки SPICE моделей транзисторов и диодов.
* Это т.н. "песочница", "лягушатник" или "черновик" для простейших схем.

*******************************************
* проверка модели биполярного транзистора *
*******************************************

* напряжение на коллекторе
VC vc 0 DC 5V

* ток базы
IB 0 vvb DC 1uA

* фиктивный источник напряжения 0В для измерения тока базы
VB vvb vb DC 0V

* транзистор
QVT vc vb 0 2N2222_LT

* SPICE модель классического импортного транзистора 2N2222
* позаимствовано из "LTSpice IV"
.model 2N2222_LT NPN(IS=1E-14 VAF=100
+   BF=200 IKF=0.3 XTB=1.5 BR=3
+   CJC=8E-12 CJE=25E-12 TR=100E-9 TF=400E-12
+   ITF=1 VTF=2 XTF=3 RB=10 RC=.3 RE=.2)
*   Vceo=30 Icrating=800m  mfg=NXP

* проверка транзистора
* -> op
* -> print v(vb)        ; напряжение на базе
* -> print i(vb)        ; ток базы
* -> print vc           ; напряжение на коллекторе
* -> print -i(vc)       ; ток коллектора
* -> print -i(vc)/i(vb) ; h21э - статический коэффициент усиления по току

*************************
* проверка модели диода *
*************************

* напряжение источника питания
VCC vcc 0 DC 10V

* токо-ограничивающий резистор
R1 vcc vd 510

* диод
D1 vd 0 NSPW500BS

* SPICE модель "стандартного" светодиода NSPW500BS
* позаимствовано из "LTSpice IV"
.model NSPW500BS D(Is=.27n Rs=5.65 N=6.79 Cjo=42p Xti=200)

* проверка диода в 

* ==============
* -> op
* -> print vd      ; падение напряжения на диоде
* -> print -i(vcc) ; ток через диод 

.end

