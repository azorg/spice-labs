* File: "lab-12.cir"
* Повышающий импульсный преобразователь напряжения (DC-DC boost converter)

* источник питания +1.5В [0.71-2.0В]
VCC vcc 0 DC 1.5V

* конденсаторы
C0 vin  0   100uF
C1 vc   vc2 2.2nF
C2 vout 0   4.7uF

* дроссель
L1 vin vl 100u

* резисторы
R0 vcc vin  1
R1 vb1 vc   1k
R2 vc  0    22k
R3 vb2 vc1  100
R4 vb2 0    10k
RL vc2 vl   1

* активная нагрузка
RN vout 0 100

* транзисторы (К-Б-Э)
QVT1 vc1 vb1 vin 2N3906
QVT2 vc2 vb2 0   2N2222

* диод 
D1 vc2 vout 1N5819

* стабилитрон
*D2 vd vout DS

* SPICE модель транзистора 2N3904 (из просторов Интернет):
.MODEL 2N3904 NPN
+  IS=6.9716e-14 BF=545.416 NF=1.09328 VAF=10
+  IKF=0.0228393 ISE=5.71808e-12 NE=1.88204 BR=4.70256
+  NR=1.3912 VAR=2.31769 IKR=0.074093 ISC=5.71808e-12
+  NC=1.36259 RB=1.733 IRB=1.12054 RBM=0.876202
+  RE=0.356192 RC=1.78096 XTB=0.1 XTI=1
+  EG=1.05 CJE=4.47982e-12 VJE=0.4 MJE=0.240345
+  TF=4e-10 XTF=1.5 VTF=1 ITF=1
+  CJC=3.76637e-12 VJC=0.4 MJC=0.241382 XCJC=0.8
+  FC=0.533333 CJS=0 VJS=0.75 MJS=0.5
+  TR=3.77901e-05 PTF=0 KF=0 AF=1

* SPICE модель транзистора 2N3906 (из просторов Интернет):
.MODEL 2N3906 PNP
+  IS=1.14615e-14 BF=535.453 NF=1.06473 VAF=10
+  IKF=0.0234918 ISE=1.33613e-13 NE=1.62939 BR=4.66099
+  NR=1.19618 VAR=2.77165 IKR=0.0740931 ISC=1.33613e-13
+  NC=1.22182 RB=0.1 IRB=1.05964 RBM=0.1
+  RE=0.0001 RC=1.39183 XTB=0.1 XTI=1
+  EG=1.05 CJE=6.03788e-12 VJE=0.4 MJE=0.272764
+  TF=4.8381e-10 XTF=1.5 VTF=1 ITF=1
+  CJC=6.18444e-12 VJC=0.4 MJC=0.234098 XCJC=0.8
+  FC=0.5415 CJS=0 VJS=0.75 MJS=0.5
+  TR=2.42096e-06 PTF=0 KF=0 AF=1

* SPICE модель классического импортного транзистора 2N2222 из datasheet:
* http://www.datasheetarchive.com/dl/Datasheet-021/DSA00361080.pdf
.model 2N2222 NPN (IS=19.34n EG=1.11 VAF=250.3 BF=163.8 ISE =174.3f
+  NE=1.647 IKF=3.0 XTB=1.5 BR=11.49 ISC=19.9f NC=1.88 IKR=10.75
+  RC=0.3567 CJC=11.02p VJC=0.3869 MJC=0.3292 FC=0.5 CJE=29.31p VJE=0.9036
+  MJE=0.4101 TR=38.32n TF=361.8p ITF=5.282 XTF=249.9 VTF=10)

* SPICE модель диода с барьером Шотки средней мощности (Imax=1A, Umax=40В)
* позаимствовано из "LTSpice IV"
.model 1N5819 D(Is=31.7u Rs=.051 N=1.373 Cjo=110p M=.35 Eg=.69 Xti=2)
*               Iave=1 Vpk=40 mfg=OnSemi type=Schottky

* SPICE модель германиевого диода 1N34 (аналог Д2Д, Д9Ж)
* найдено где-то в сети Интернет
.model 1N34 D(Is=100p Rs=84m N=2.19 Tt=144n Cjo=4.82p M=.333
+             Vj=0.75 Eg=0.67 Bv=60 Ibv=15u)

* SPICE модель абстрактного стабилитрона (импровизация):
.model DS D(Bv=5.6 Ibv=5m Is=2.52n Rs=.568 N=1.752 Cjo=4p M=.4 tt=20n)

* температурный режим
.options TEMP=25

* моделирование переходного процесса
* шаг моделирования - 1 мкс
* время моделирования - 0.1 с
.tran 0.1u 10m

.end

