* Лабораторная работа №3
* ----------------------
* Файл: "lab-3_1.cir"
* Измерение входных вольт-амперных характеристик (ВАХ) 
* SPICE модели биполярного транзистора

* напряжение на коллекторах транзисторов
VC1 vc1 0 DC 0V
VC2 vc2 0 DC 0.5V
VC3 vc3 0 DC 0.7V
VC4 vc4 0 DC 2V
VC5 vc5 0 DC 15V

* напряжение на базах транзисторов
VB vb 0 DC 0.5V

* фиктивные источники нулевого напряжения для измерения токов баз
VB1 vb1 vb DC 0V
VB2 vb2 vb DC 0V
VB3 vb3 vb DC 0V
VB4 vb4 vb DC 0V
VB5 vb5 vb DC 0V

* четыре одинаковых n-p-n транзисторы с разными напряжениями на коллекторах
QVT1 vc1 vb1 0 KT315B
QVT2 vc2 vb2 0 KT315B
QVT3 vc3 vb3 0 KT315B
QVT4 vc4 vb4 0 KT315B
QVT5 vc5 vb5 0 KT315B

* SPICE модель классического советского транзистора КТ315Б (h21э=100)
.model KT315B NPN(Is=14.34f Xti=3 Eg=1.11 Vaf=125 Bf=124 Ise=157.3f
+  Ne=1.558 Ikf=.2999 Xtb=1.5 Br=1 Isc=15.86f Nc=1.022
+  Ikr=3.163 Rb=15 Rc=3.748 Cjc=8.988p Mjc=.33 Vjc=.75 Fc=.5 Cje=18.5p
+  Mje=.33 Vje=.75 Tr=301.4n Tf=321.4p Itf=1 Xtf=2 Vtf=60)

* температурный режим
.options TEMP=25

* DC анализ при различном напряжении на базах (0...1В)
.dc vb 0V 1V 0.1mV

* Гграфики зависимости тока базы от напряжения на базе
* -> run
* -> plot i(vb1) i(vb2) i(vb3) i(vb4) i(vb5)

.end

