* File: "lab-3_3.cir"
* Анализ зависимости тока коллектора от тока базы биполярного транзистора

* источники напряжений для коллекторов транзисторов
VC1 0 vc1 DC -1V
VC2 0 vc2 DC -9V
VC3 0 vc3 DC -20V

* заданный ток базы транзисторов
IB 0 vb DC 10uA
VB vb 0 DC 0V

* трансформаторы тока для размножения заданного тока по базам транзисторов
F1 0 vb1 vb 1 m=1
F2 0 vb2 vb 1 m=1
F3 0 vb3 vb 1 m=1

* идентичные n-p-n транзисторы с разными напряжениями на коллекторах
QVT1 vc1 vb1 0 KT315B
QVT2 vc2 vb2 0 KT315B
QVT3 vc3 vb3 0 KT315B

* SPICE модель классического советского транзистора КТ315Б (h21э=100)
.model KT315B NPN(Is=14.34f Xti=3 Eg=1.11 Vaf=125 Bf=124 Ise=157.3f
+  Ne=1.558 Ikf=.2999 Xtb=1.5 Br=1 Isc=15.86f Nc=1.022
+  Ikr=3.163 Rb=15 Rc=3.748 Cjc=8.988p Mjc=.33 Vjc=.75 Fc=.5 Cje=18.5p
+  Mje=.33 Vje=.75 Tr=301.4n Tf=321.4p Itf=1 Xtf=2 Vtf=60)

* температурный режим
.options TEMP=27

* DC анализ при различном токе баз (0...1mA)
.dc ib 0A 1mA 0.1uA

* Графики зависимости тока коллектора от тока баз
* -> run
* -> plot i(vc1) i(vc2) i(vc3)

.end

