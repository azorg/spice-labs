* File: "lab-1-simple.cir"
* Изучение усилителя переменного тока на биполярной транзисторе с
* по схеме ОЭ и обратной последовательной отрицательной связью по постоянному
* и переменному току.

* конденсаторы
CIN vin vb 10uF
COUT vc vout 100uF
CE 0 vce 33uF  
CVCC Vccc 0 1000uF  

* резисторы
R1 vb Vccc 47k
R2 vb 0 10k
R3 vc Vccc 3.3k
R4 ve vce 100
R5 0 vce 1k
R6 VCC Vccc 100

* внутреннее сопротивление источника
RIN vsin vin 1k

* сопротивление нагрузки
RL 0 vout 3.3k

* источник питания +9В
VCC vcc 0 DC 9V

* источник сигнала
VSIN vsin 0 dc 0 ac 1mV sin(0 1mV 1kHz)

* n-p-n транзистор(ы) (C-B-E)
QVT1 vc vb ve 2N2222

* SPICE модель классического импортного транзистора 2N2222 из datasheet:
* http://www.datasheetarchive.com/dl/Datasheet-021/DSA00361080.pdf
.model 2N2222 NPN (IS=19.34n EG=1.11 VAF=250.3 BF=163.8 ISE =174.3f
+  NE=1.647 IKF=3.0 XTB=1.5 BR=11.49 ISC=19.9f NC=1.88 IKR=10.75
+  RC=0.3567 CJC=11.02p VJC=0.3869 MJC=0.3292 FC=0.5 CJE=29.31p VJE=0.9036
+  MJE=0.4101 TR=38.32n TF=361.8p ITF=5.282 XTF=249.9 VTF=10)

* температурный режим
.options TEMP=25

* моделирование переходного процесса
* шаг моделирования - 1 мкс
* время моделирования - 10 мс
.tran 1u 10m

* AC анализ слабых сигналов при снятии АЧХ/ФЧХ
*.ac oct 3000 1Hz 100MegHz

* контроль рабочей точки по постоянному току:
* -> op
* -> print v(vb) v(vc) v(ve) v(ve2)

* симуляция переходного процесса
* (анализ переменных напряжений на входе и выходах
* -> run
* -> plot v(vsin) v(vout)

* снятие АЧХ/ФЧХ (1Гц...100MHz)
* -> ac oct 3000 1Hz 100MegHz
* -> plot db(ac.v(vout)/1mV)
* -> plot ph(ac.v(vout))*360/(2*pi)

.end

